`timescale 1ns / 1ps

module mux16bit(
input [15:0] in0,
input [15:0] in1,
input sel,
output wire [15:0] out
);


endmodule
