module train(
    input rx,
    output tx,
    output [7:0] led
);

endmodule